module dm74ls283_quad_adder_tb();

input reg [1:4] a, // input b
input reg [1:4] b, // input a
input reg c0, // carry in
output reg [1:4] s1, // sum
output wire c4 // carry out

// todo

endmodule