`default_nettype none
module ram(
    input wire [7:0] dipswitch_data,
    input wire [3:0] dipswitch_addr,
    input wire [7:0] bus_data,
    input wire addr_button,
    input wire data_button,
    input wire write_enable,
    input wire output_enable,
    input wire control_signal,
    input wire load_addr_reg,
    input wire clear_addr_reg,
    input wire enable_addr_reg,
    input wire clk
    output wire bus_out
);

  wire [3:0] mem_low, mem_high;
  wire write_mode;
  wire run_mode;
  wire address;

  sn74ls159 mux1 (
      .a(dipswitch_data[3:0]),
      .b(bus_data[3:0]),
      .select(data_button),
      .strobe(0),  // output always on
      .y(mem_low)
  );

  sn74ls159 mux2 (
      .a(dipswitch_data[7:4]),
      .b(bus_data[7:4]),
      .select(data_button),
      .strobe(0),  // output always on
      .y(mem_high)
  );

  sn74ls159 mux3 (
      .a(run_mode),
      .b(addr_button),
      .select(data_button),
      .strobe(0),  // output always on
      .y(write_mode)
  );

mar addr_reg(
    .dipswitch_input(dipswitch_addr),
    .button_select(addr_button),
    .clk(clk)
    .bus(bus_data[3:0]),
    .load(load_addr_reg),
    .clear(clear_addr_reg),
    .enable(enable_addr_reg),
    .mar_out(address)
);

assign internal_data = {~mem_high, ~mem_low};
assign run_mode = ~(clk & control_signal);
memory mem(

    .data(internal_data),
    .write_enable(write_mode),
    .enable(0),
    .address(address),
    .bus_out(bus_out)

);
endmodule