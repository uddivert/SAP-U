module dm74ls283_quad_adder(
    input wire [1:4] a, // input b
    input wire [1:4] b, // input a
    input wire c0, // carry in
    output wire [1:4] s1, // sum
    output reg c4 // carry out
);

// todo

endmodule